library verilog;
use verilog.vl_types.all;
entity decoder_top_tb is
    generic(
        PERIOD          : integer := 10;
        CW_W            : integer := 16
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of PERIOD : constant is 1;
    attribute mti_svvh_generic_type of CW_W : constant is 1;
end decoder_top_tb;
